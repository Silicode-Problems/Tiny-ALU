module tinyalu(
    reset,
    op_code,
    A,
    B,
    out
);
 // Your code here   
endmodule 
